library verilog;
use verilog.vl_types.all;
entity nios2_tb is
end nios2_tb;
